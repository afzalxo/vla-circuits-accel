`timescale 1ns / 1ps

module conv_accelerator #(
    parameter IC_PAR = 16,
    parameter OC_PAR = 16,
    parameter PP_PAR = 8,
    parameter DATA_WIDTH = 8,
    parameter MAX_IMG_WIDTH = 128
)(
    input wire clk,
    input wire rst_n,
    input wire start,
    
    input wire [15:0] img_width_strips,
    input wire [15:0] img_height,
    
    input wire signed [OC_PAR-1:0][IC_PAR-1:0][DATA_WIDTH-1:0] weights,
    
    input wire signed [PP_PAR-1:0][IC_PAR-1:0][DATA_WIDTH-1:0] din_data,
    input wire din_valid,
    output wire din_ready,
    
    output wire signed [PP_PAR-1:0][OC_PAR-1:0][27:0] dout_data,
    output wire dout_valid,
    output wire done
);

    wire lb_shift_en, seq_load, cu_en, cu_clear;
    wire [1:0] k_x, k_y;
    wire [15:0] col_idx, row_idx;
    
    wire signed [PP_PAR-1:0][IC_PAR-1:0][DATA_WIDTH-1:0] row_0, row_1, row_2;
    wire signed [PP_PAR-1:0][IC_PAR-1:0][DATA_WIDTH-1:0] seq_out;
    
    // NEW: Wire for valid out (unused but good for debug)
    wire cu_valid_out;

    conv_controller #(
        .MAX_IMG_WIDTH(MAX_IMG_WIDTH), .PP_PAR(PP_PAR)
    ) ctrl (
        .clk(clk), .rst_n(rst_n), .start(start),
        .img_width_strips(img_width_strips), .img_height(img_height),
        .din_valid(din_valid), .din_ready(din_ready),
        .lb_shift_en(lb_shift_en), .seq_load(seq_load),
        .k_x(k_x), .k_y(k_y),
        .cu_en(cu_en), .cu_clear(cu_clear),
        .col_idx(col_idx), .row_idx(row_idx),
        .dout_valid(dout_valid), .done(done)
    );

    line_buffer #(
        .IC_PAR(IC_PAR), .PP_PAR(PP_PAR), .DATA_WIDTH(DATA_WIDTH), .MAX_IMG_WIDTH(MAX_IMG_WIDTH)
    ) lb (
        .clk(clk), .rst_n(rst_n), .shift_en(lb_shift_en), 
        .img_width_strips(img_width_strips),
        .data_in(din_data),
        .row_0(row_0), .row_1(row_1), .row_2(row_2)
    );

    window_sequencer #(
        .IC_PAR(IC_PAR), .PP_PAR(PP_PAR), .DATA_WIDTH(DATA_WIDTH)
    ) seq (
        .clk(clk), .rst_n(rst_n),
        .kernel_y(k_y), .kernel_x(k_x), .load_new_data(seq_load),
        .col_idx(col_idx), .img_width_strips(img_width_strips),
        .row_idx(row_idx), .img_height(img_height),
        .lb_row_0(row_0), .lb_row_1(row_1), .lb_row_2(row_2),
        .pixels_out(seq_out)
    );

    vector_compute_unit #(
        .IC_PAR(IC_PAR), .OC_PAR(OC_PAR), .PP_PAR(PP_PAR), .DATA_WIDTH(DATA_WIDTH)
    ) cu (
        .clk(clk), .rst_n(rst_n), .en(cu_en), .clear_acc(cu_clear),
        .valid_in(cu_en),
        .img_vector_in(seq_out),
        .weights_in(weights),
        .img_vector_out(dout_data),
        .valid_out(cu_valid_out)
    );

endmodule
