�      �=kw�6����
4MZ:ud�~�vݻ��ĺ�%�$7=��GKK�Ř"�$�Ǿ~���A$HK��v���$��`03����0��W��O�Z|�䑟:<[[����i����؛��O�M۩ۛ���擺��������3�7"�;���W����?��K�Mi<t}J� &kĞ�ϞM��Jr�A���xfn�NiǍ��������!�#��f5���dp��Bݛg+����	��"����/��dJq�^��:�7w��ě^n�Q2�I����J�	�.'%Í�`p��ވW���"z�j"�J�1�'�8Р�5���[��F����5w�����	(�ԍ����C��Lc�Qx�U���0����3V�@N� Ho�:8j���n��I�u�t;X{����#@�7�^־���������^%=\}CG�p�i��;oX�V $:�#�M���IHfs?��UA��H�%إ��?�����i�)��a��F���}���]��8h7�c��lmz��9:���a�:��Ο�ҥS������[�z�i+��-���:���n���F����L��Ċ� A��\��W�Agތ�4�eծ����O�,����&F$��앉�rA/�����7&�7�|�r��'�`W�L�	6��u�$1�J�0T1�`.g���)W�!_���R�P#�iN�j�U��2T+t`��4׀#B����{@���O�	r\�8�P@�S�5������NM;��d �M>H�l?5����5+4-_?mr�ԣ>唤>
�����5�A��
��N�_�&v��ɯ�n���8"ېV��ԩ�w�9� �o��1��� $�N_����C(7,k:�ʵUix�)#������7������b�(�ȷ�^�pc�A<gzu����Vs���V��4r��+h�V����٧�ү�>�e�Ly�
�u���U�������k�5��n��:�>���9'S�JY����럹H�8�X�<ߏ���'ߛĢ���p����J1��(���q��~]�Z�����$�]�&]`o��*���E�W�F�-[x`g�{�|pM
k ����a-TL�Yi��R�Eɭ�;Kn�O�fcI��ܦS�,4IFk�DκA�89�c��Σ��U0q�� ��*���C��6pș�{M�9�px:�Y�B�v6��9��/��[.x*J��6��'�}�M���=�k�c/'z��U����^�hIǩH��ȏ��nj�W`]]�
�_w� ��������/+�닯�����R��P�J�@�Q�=g�[���d6k���#�'�R��6�QMnr 7��+QA>Ur�t6BDu��w?#��PR)����	�z1�>��@�|,� !>Ȩ§
��:�"�0b٧������D-���}�;Ћ� 2ӝZn�?����9/|�Y
emĥ��|�L���n�(Ir%U�l)�y�F脹�{�n�Rq��UW(z��� e2U�n�H́+�^��.�x�%3^>��$�XH͙a��"�q�z
���n�4�؇ �KoH�����@���7f�@����#/0X2���P�΅�(�_N����jxA�*y�B�<�
S_�S�䔦����W��|L3����)�vy�9��B���f����Q������>>K�'�uN����S���$��=eu��T$�lg2��pK�'��!,R�R���ÈN)����>�_ ��^�P&1��Ry��T�-)�{+�,R�6��#���H>
���Y6�qK��"a�
G�7"NVʕ���1��,_�@��x�ͳ�;��Im��:�������§:����i���/{����_�u�k�חx*��(�~��Eb��U�����f�j��d��֧%�i�XH��� T�3>�ט�u���g�a�L_x��?��af,���
)E�5�'w�%�u�������U�4���<B1>T�w�o� �P��We�q�qL�b����y�_'�5AT�j�W��������D�s�k�,�nY�`�:9��p���w?��l���1��D�Yr��/���d��#�6߷z�f����PߟP��'�?b���:,��2;GP�MX�;�4C�Y�w?q �Spd�W��9/�j�)uvZgꜴ����
��;�o	�X=o:�]�ڰpߊ�*	���W�'�� �-�%J���������ɪa�{杓��ͨ�P�i#b�oB�������'�q�7����*����إ5N._+�^YNK����Y2Q��8 '��^�X��,�4�C�atWN��M����G��پT��y2�_��x�w�sL�%�dB�'n j�y9Z���|Ux�^?�^m���_����uS��_��u�")NCJ��K�q�}��C�!^��&�@a����	XF<)�~Ias�1��������9�	7�-�%�c��˨���2L��BB���.c .ү�hө��V�)�S���h�Cn@o��(��M,�uAAi��('�b�\{�of���i�bU���5����1�6������1�#  �� �3�V�C�Ä� ��J#�/A[^_�zr�����-M[M��l9������9Fh�����)q����>�1��W��lc�
p�f�Wj�1{��!ȅa�ߑ)�@!a��9@������YVaZ&[tZm�,�bX(��^�-W*��e��_Z6��e��e��_�V�}�G����֦�p�@(���r������{k{s���κ�����O��/I���W�E��_l������7l�O1���Ϙ�8u��;�*Y���g��Jv��w�t�r/BU����'�� )΄uCc0C��8���L��I3��7��fV�?���p�ny#�^�H�E�;�~�s�>y�j�n��[� S)>���l:�������;�Wj���DN�l�)�2��� @�)=Z� ��٫�Pgub��I	������?�wg��!�̹>
A�SZl��2e�(�����Q�D���^.�K��߳�"�){����T(sD�.z�#fH7�»Y3 ��D��)���T�����$M���t0�g��1�z4f�>@�h>⬾#���谰����t�3�϶��v���6�6?27c�ć�\rޅ��X�5������D�מ��s�f0��J�]�dr�G�h!�pc�?

���^�ǖ"ɡf��Jk���ҥt��.Tʣ�1���#
FC�/y4��\̅� &S�tAI}�t=ߤ�p
�a$�y���X�Ǌ���N�������9���>��9g0���:�����,�ҕX{U�l&�*��D^�m±�G��I#mC^8�n����<<Ǎ}0[a�wHc����T��?`x��=��)'{T�G�.)�u���
��Z�D,�-�ǧG�~��9�~�-%d �a�%wr��8�3�mQ�h[Q���S��L��hR3����G�hH��*3��(�����}z�=lP�z�%�m�8�7^L�ϣϝ��Ҷ��?$C(���H���ʍQ��vM]HK�ڔ���&�%*���U�N�(w�a�Y����}jk��!�)�P��<�'����ܮs��q�6ס��������/�T��E�X*�S^��>��/��K�}e_�{�MNp�%��%%1���^��C�z�i>�7�>�E�y>���-Q>�~���F�w��o?h#z{~&:�׷^"~���_,�'v��\�<�����0}����m�a��e��M��i�v6�EtI�k`��]�F#u�gj���^����=��`a+|�l�����{�ԧƑn�VV��������BpxXP� ֱP5�8��
�����*R���_���Ӛ�'K�0�V4HKrĊp�M��@�b�5�v�(P]q}�M4.�(�������\��R�;_�N&�@#��K�yB�9 I��Z��q�J)����J,���R_�J���P���%��܇5�0�g	T����������t���o�_����S��k��{�@z5��Z���dV���|]��.K,T�C��pݮ�s�X?��e\舝��7i�1+��NZ�z��Һ��7��և�6���^�}L���7Њ��o����\f�$�]Pp.����@3�cz�Dq̦�<t�rS����G��:"	�4�g���ٌ8��qH�0���q��m5�e�{���*?zO�}��k�ae�7r�Tk�ڽ~��o5��N;�]��2h�ф��z�U��Q�0X�b�����j����BcEK{��
�U�%�X�Q4UE)gd/���t���d<>�t�B-�� Z���706�(��&?O���4�~kC*.��po�A^9Q��Iβ�mj)�e'�
���찗��ܭ��>NJ�V�3�"��%,�;�����o������}�ɜy{�_����]�)sT�#��dc���n�ȿ���ܯE���2�����ů�J�$fM5o�����o���0RɒoE�)uF�kj*hD��g��QFEZ;W�;W����<�)lz�
�S��D�-Z��*��d��z�v�3kz�|U
0E�U��MorE-��j2�����^����'7n�Ն�5���2.��x��7PO�$����\�B��p*��z�8[�1�c*	'��֩�k��a�\6�خ+�i\�>�^��������(�O}��(
����(#�U<��Ɠ�̱)��7促n��f︹���n0�'���/��(�p�bJ��8���fD{�?F�y&�e~+f��a�{;���s~�L��x���)h��Vu�TJt�����t�\f�=��4á�B�!�Ij�
�l��|
���YB�1��y�	b��$��p��G��}s�^����E��EZ�O��U�N�3dySq��G�oF��v�R�t��_̖��C�RA�����S���	z��Q�6���;.�b*d�	�,���T'Pr��C�U?���D����@�F�^97{6hs��xGf���j��C�%�P9�;�����l��3'L2OQ�ʒ%f|�k}�MH�hVv�#�8������U�y1fY��fak{Yǈo+�����l�E�Շ:�/���]}n�j:�����A��)���A5L;���� פo?�� �RW5r`�}Xnhi�QZ%u�BeV�'σ����;�e �=}���<��<��D;�,�Tm�]������P�^��K��lU�XT�>v��zB�Azx����}�N��0	�;�/@%i/����aͿ���7eO�N_y��=Fxj��Q�:��� ����6Yj:����{�]դ	^������''�Ĉq�}����
�4�bc���]�,��va�c
���^�mb�����ۏx�X�K ^_����~�!���O����䅸�/��˅ȵG�RV�dکBp�Js���R~�r��r�
��d|��.�����b��\����H�uw���*�c�%ATw��?��/���?��b��N���2Fx���Y����fe�"M�jÏC��t��x�7ܘ*ǲ|4p�h\��h]z�Uq�֙�}P�_Ǩ�rw"����9ٿǜ��;'������`��B��ƌY��	|�/��{��<�kom�;�S�������__�/���F��?��&�%��H����N�آj>��H�p�F>���+*�CΟp�������)�f�^~~��1���f��Ԧ�䅲T(Z�n���,��	�D���������4�⊳�'-�r��F�I/w��Dj?�%M�HC3̵*#4Y(�%��e�c~+~h8#���ol��+�6õN�Ņ(pi�w���a��"��ݟݫ�F&Q�|�n�e��*�4���:�������a�����d��G��@�@� ���F������P���5.��7u���f����[�e5W.vU�ѿ�@�(� J�B(��lK�}����` n��Q:T�T>bɥ��m�j&��S)&f���N�bbP-�4Ȳ!M�Jwě�M�7�T�O�����ͣ�f���_4�ށ�3ja@���̓�M����i2��C��Li"���g,�Ot��zC���N�č�Ș��X�7Co LPѵӓ���cVZt`�ɒ'�pi����Y���c�!��Da��,=u���pҦ��
�l��~LO~��hl���C�;?�x�Ӟ�-xt�w��D�|2������i�%o0�Jfe�T��>;yY�`ҁ!�P��E� l|t)�1-�`#�����`�j��ɲ�Q�|��Ƣ^Hmxki�3�l��Bc�~��/D�26(Ms���+z6	NXͷ�w{���6r��o�)x��Y�.e�q�E~ :+�"��$Bd���T���ξ8�")�v��<lr�;;ܝ���.	(	b4�����b"Gxi��94�&��w�P�{]iy��o��ZÒ�0���Ny��u*�!�G�wzxr�� '���ȧ??@E^ G
u	��d���LeG�+3���;�B��N��^IQ�*�D@�"[d�h�,��~�Y�$��{rzdX�jl܁ude�l��rȾ"�0G0ܱ0�"���1�E���IT��_&�e��@�bX�O�%K:dL��P?���AG�7|ju{_�BU���`Nd掮���׽4����0�8��i���jp\�E�quj�-4A`󄟩0�G5�=,���J�?���H��C�9�����_-!D�GI�����y�w#�D�X���}[1Zؘ��-��w�_�M~���/'��u-�����D�|Qcm*�����/�@��E#�M1@ pR�T��t?-�c��-I�H@%�d���`�_��"�7�[y���W�o�nRB�휞�
L�'���ҁ�-��-Q/�6wd�'&/��w�{镠ۋ�k�(� &;'�R�`į�K�dLZ;@J���V��l�I�KR.:f�|
����v��3���k�[_A�#a�]τ���1R,RNː��Z�k< �$�,�@ze��Ū�-����62"�ۈӃnt�9��^�_�,��y9�{�Gj��lğ��l��SzJ���'�j���B�l��o����������ێa9� �<8�|�[gc�l�O]sk4��H���
��5(�ip�x:�yxpҽ<��EU�݈>Mf~�0v�����K6�1`�b�}.k腍�ηr����(����K����d���?lW�����5ֱ�=������T�Nno�(��h��W�j�e��F�|-��p�� K35���@4e�}�q4����QHX���.�}\��
j�����IURfc4�K����?�
9�y���p���zB�'T=~��]O?���GG���-/ijf�n�G��T63�[���B�6��M�G�Qo������~<���)@�P�쨛/��}���=��QqjRc�FV�(�У	k'�hhx4x |uL١�٨��^A�����l����euc�Vkf��w��~ŷG�й{��-a/���}�8�q��T�`����^t�鼊�zo�&s��1a�$����7� Ĳ��M���1��HO���Դm�ڥ'H�lH�Rh,��a��6���,����l�dl}�K�a�on눯u��|{��b_���B�B�Ԯ��+L����S�}�'+ԟ��'v��Q�tD3eY)7ʺB�`:V���~�2����WZ��������}����#���_�9<C��yC��}ؚ���ݲ�����15�FB�-G(�&�i�<�=U�O0�dn�,sgSb׸w�e�X�R��{�j\����ibט��	bh�:aE%,{��,�Ь�C���.�j�.'M������*żJ\5y9���=Ţ4Ȣ�`���c��c�}cf�«��a�F��s�mh#���z|5�y:��N7w(U|���*�6]b8jg�F;��-����Ӕ2n��c��@h��B�bm�����!���Qm��*���j��m����iU��Ǡ"�����*V�`�� 憲�7�h�n9S�pQPK@vNW�@��k�hr�,ȸ����2�f@���@ڒJ�,����h����Ҫ4��! ��~\F��a=�R�l�2��V��z��n�P�߉�;�(�2o@~��2�U��j��mR����Y��:����09�ɩ?y�3�<�����q��Z��0&��j�lI׭\Tb��NlxI���%U]<֭��iظ�� (��9���[rM[��o�\��+���Z�0��N�N���S?����n�
�4qF�ht_h�d��	E�@�X��(�3��p<gX�Qu������3+��������8�p�(t0^Xa�p���#�h�f�s`����ٽWe���ڧA���8▒ftί��].P�5h���HOWv�ˁBzq��)�屖�50y��ϓ�1��x��4R�`�1�g0v������⯮@X׺�ɗ�2��e�P�`.z��H|�n �V�$U^�~४�=��M��
��}V��a�d$��ߌ�_�~+��0!���OvVɵF45s���� �mZ�&f��>s��яF�f�z��V�V�67�;Dm5DǓ���&73g��Ï3{�tk�@kٟhrf����������ܝO��W0��pƁ����{�Fʮwzqrzyr��`3�X'���r)E��~:�C�!�3��=���'q�l9��r
�!yB%Or�z$����)|�~��Ҭ�KTȺ�G5>jm���occ�+���܃����t�	Q�5�k��6=�x�_n1a�VE�N�[�WY8{�[�$�/��F��4ںVXt|b7��l��%\�U��k�G�#V�cRs�sW�Q��q�m���\���T��Ǡ\�o�5�u@e�������r�h0��X9�/CF�V�7��x7�U����;�2����?��L��j�}�*9��8S�>9�k��O�R�<%�(��S%����SoN~�t��S�xm��cPY����T�?P�*��f��w�{"(�B@)7+/������3���gz��!܎� g�5�	F��P�L���
�J��T=5�����b���6�����g���I+���A�����������y'g��  �5���}o9�����M��.� �P�ʔ(��p���d:#�*�
�h��m�Cf��;:i=���!�@�%�
�M��4Crc�>ҫ4��]��U��R
�nt
�0d�A����<�_E����� �w��F�Q)���M�Q�)2�!ۍ�A�9�:��Sw r���å� �p��/����e�[�����E�8���N�Y��w� �u�����;?"�Oyt%8Jj��ͦ�/��`#��dO���D%����[�DCэ`�L$������:�.��1(��|���r�΀�A1�T��bE��5(��Z)�hw�6���K��_T�r��)��v�Fh:=�53��ԴA�
M6�<j��<�JE��(JE��93d��orao���˻[��W�YN�鬜�8o�r�[�!7��l�vݔa����Cy���z��²� VQMm?ͳ7}z�I������MD�$���¨3��Ʀ�j��^;N���ͭ�(��F��9�@(���}�t�K�\��z<��#/{�_�f��
�� ]~��:�쫯 r��LZ��<؆����/|�Y����|Q��W
�e,ع�w�-��#���|$wͪ�-��cX�{�/�3ް_0���NQš�r�N|�:[ T|!� ��ܐ,㭢�i���m ^�g�L�']}��8��{}p�9x%��e���E��R�_N�n�����6E%9D��r:�o߫0C<�c8�b��� �Iκ�D�&�.�_?��7#w>l�E&.�BfTTQEUTQEUTQEUTQEUTQEUTQEUTQEUTQE��O�P] �  